`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:08:07 03/16/2016 
// Design Name: 
// Module Name:    data_mem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`define idle	1'b0
`define exec	1'b1
// instruction 
`define NOP	5'b00000
`define HALT	5'b00001
`define LOAD	5'b00010
`define STORE	5'b00011
`define SLL	5'b00100
`define SLA	5'b00101
`define SRL	5'b00110
`define SRA	5'b00111
`define ADD	5'b01000
`define ADDI	5'b01001
`define SUB	5'b01010
`define SUBI	5'b01011
`define CMP	5'b01100
`define AND	5'b01101
`define OR	5'b01110
`define XOR	5'b01111
`define LDIH	5'b10000
`define ADDC	5'b10001
`define SUBC	5'b10010
`define JUMP	5'b11000
`define JMPR	5'b11001
`define BZ	5'b11010
`define BNZ	5'b11011
`define BN	5'b11100
`define BNN	5'b11101
`define BC	5'b11110
`define BNC	5'b11111
//register 
`define gr0	3'b000
`define gr1	3'b001
`define gr2	3'b010
`define gr3	3'b011
`define gr4	3'b100
`define gr5	3'b101
`define gr6	3'b110
`define gr7	3'b111

module data_mem(reset,mem_clk,dwe,addr,wdata,rdata,tocache);
input reset,mem_clk, dwe;
input [15:0] addr;
input [15:0] wdata;
output reg[15:0] rdata;
output reg[63:0] tocache;
reg [15:0] d_mem[2048:0];

always @(posedge mem_clk or posedge reset)
begin
  if(reset)
  begin
  rdata <= 0;
  tocache <= 0;
  //������� ��С������data
  /*d_mem[0] <= 16'h0000;
  d_mem[1] <= 16'h0020;
  d_mem[2] <= 16'h0018;//*/
  
  //ð������data
  /*d_mem[0] <= 16'h000a;
  d_mem[1] <= 16'h0004;
  d_mem[2] <= 16'h0005;
  d_mem[3] <= 16'h2369;
  d_mem[4] <= 16'h69c3;
  d_mem[5] <= 16'h0060;
  d_mem[6] <= 16'h0fff;
  d_mem[7] <= 16'h5555;
  d_mem[8] <= 16'h6152;
  d_mem[9] <= 16'h1057;
  d_mem[10] <= 16'h2895;//*/
  
  //sort
  /*d_mem[0] <= 16'h000a;
  d_mem[1] <= 16'h0009;
  d_mem[2] <= 16'h0006;
  d_mem[3] <= 16'h0005;
  d_mem[4] <= 16'h0001;
  d_mem[5] <= 16'h0004;
  d_mem[6] <= 16'h0003;
  d_mem[7] <= 16'h0011;//*/
  //cache
  d_mem[0] <= 1024;
d_mem[1] <= 13962;
d_mem[2] <= 6923;
d_mem[3] <= 10905;
d_mem[4] <= 22204;
d_mem[5] <= 21127;
d_mem[6] <= 7322;
d_mem[7] <= 18464;
d_mem[8] <= 6849;
d_mem[9] <= 604;
d_mem[10] <= 23895;
d_mem[11] <= 320;
d_mem[12] <= 16557;
d_mem[13] <= 22383;
d_mem[14] <= 8835;
d_mem[15] <= 8972;
d_mem[16] <= 4911;
d_mem[17] <= 22509;
d_mem[18] <= 9623;
d_mem[19] <= 15522;
d_mem[20] <= 16988;
d_mem[21] <= 24253;
d_mem[22] <= 15927;
d_mem[23] <= 23265;
d_mem[24] <= 25939;
d_mem[25] <= 11430;
d_mem[26] <= 341;
d_mem[27] <= 3939;
d_mem[28] <= 7742;
d_mem[29] <= 2510;
d_mem[30] <= 8982;
d_mem[31] <= 16688;
d_mem[32] <= 393;
d_mem[33] <= 25786;
d_mem[34] <= 24221;
d_mem[35] <= 9544;
d_mem[36] <= 11209;
d_mem[37] <= 13810;
d_mem[38] <= 7585;
d_mem[39] <= 2116;
d_mem[40] <= 19509;
d_mem[41] <= 3009;
d_mem[42] <= 23906;
d_mem[43] <= 11367;
d_mem[44] <= 20833;
d_mem[45] <= 2447;
d_mem[46] <= 7154;
d_mem[47] <= 8777;
d_mem[48] <= 18537;
d_mem[49] <= 20796;
d_mem[50] <= 12271;
d_mem[51] <= 5347;
d_mem[52] <= 18658;
d_mem[53] <= 25918;
d_mem[54] <= 252;
d_mem[55] <= 7154;
d_mem[56] <= 20218;
d_mem[57] <= 25918;
d_mem[58] <= 2805;
d_mem[59] <= 5478;
d_mem[60] <= 12255;
d_mem[61] <= 17471;
d_mem[62] <= 23775;
d_mem[63] <= 3677;
d_mem[64] <= 4086;
d_mem[65] <= 1050;
d_mem[66] <= 12854;
d_mem[67] <= 13925;
d_mem[68] <= 25393;
d_mem[69] <= 7784;
d_mem[70] <= 21626;
d_mem[71] <= 17634;
d_mem[72] <= 23228;
d_mem[73] <= 7737;
d_mem[74] <= 7905;
d_mem[75] <= 9838;
d_mem[76] <= 14792;
d_mem[77] <= 23901;
d_mem[78] <= 25445;
d_mem[79] <= 9192;
d_mem[80] <= 9198;
d_mem[81] <= 23354;
d_mem[82] <= 14965;
d_mem[83] <= 12234;
d_mem[84] <= 8425;
d_mem[85] <= 15785;
d_mem[86] <= 13883;
d_mem[87] <= 24100;
d_mem[88] <= 16205;
d_mem[89] <= 12113;
d_mem[90] <= 13741;
d_mem[91] <= 24137;
d_mem[92] <= 1507;
d_mem[93] <= 19630;
d_mem[94] <= 13510;
d_mem[95] <= 4832;
d_mem[96] <= 7653;
d_mem[97] <= 18012;
d_mem[98] <= 2479;
d_mem[99] <= 4338;
d_mem[100] <= 21048;
d_mem[101] <= 16788;
d_mem[102] <= 9985;
d_mem[103] <= 19131;
d_mem[104] <= 777;
d_mem[105] <= 4916;
d_mem[106] <= 13846;
d_mem[107] <= 12176;
d_mem[108] <= 12334;
d_mem[109] <= 17702;
d_mem[110] <= 7601;
d_mem[111] <= 20344;
d_mem[112] <= 9712;
d_mem[113] <= 24468;
d_mem[114] <= 25366;
d_mem[115] <= 472;
d_mem[116] <= 13594;
d_mem[117] <= 10274;
d_mem[118] <= 9297;
d_mem[119] <= 26159;
d_mem[120] <= 20203;
d_mem[121] <= 8683;
d_mem[122] <= 12717;
d_mem[123] <= 23985;
d_mem[124] <= 12355;
d_mem[125] <= 2432;
d_mem[126] <= 78;
d_mem[127] <= 3593;
d_mem[128] <= 2017;
d_mem[129] <= 16063;
d_mem[130] <= 13909;
d_mem[131] <= 2216;
d_mem[132] <= 3172;
d_mem[133] <= 1780;
d_mem[134] <= 16494;
d_mem[135] <= 3025;
d_mem[136] <= 5442;
d_mem[137] <= 2946;
d_mem[138] <= 914;
d_mem[139] <= 8877;
d_mem[140] <= 562;
d_mem[141] <= 13515;
d_mem[142] <= 3803;
d_mem[143] <= 4622;
d_mem[144] <= 998;
d_mem[145] <= 7616;
d_mem[146] <= 10353;
d_mem[147] <= 22377;
d_mem[148] <= 2316;
d_mem[149] <= 11041;
d_mem[150] <= 22251;
d_mem[151] <= 4885;
d_mem[152] <= 24615;
d_mem[153] <= 14408;
d_mem[154] <= 8441;
d_mem[155] <= 21962;
d_mem[156] <= 16846;
d_mem[157] <= 14419;
d_mem[158] <= 18317;
d_mem[159] <= 8362;
d_mem[160] <= 10621;
d_mem[161] <= 2600;
d_mem[162] <= 18275;
d_mem[163] <= 3067;
d_mem[164] <= 22666;
d_mem[165] <= 25261;
d_mem[166] <= 10227;
d_mem[167] <= 20255;
d_mem[168] <= 9528;
d_mem[169] <= 5531;
d_mem[170] <= 12785;
d_mem[171] <= 5321;
d_mem[172] <= 9187;
d_mem[173] <= 17313;
d_mem[174] <= 4465;
d_mem[175] <= 13631;
d_mem[176] <= 17145;
d_mem[177] <= 1292;
d_mem[178] <= 24100;
d_mem[179] <= 4911;
d_mem[180] <= 14892;
d_mem[181] <= 19000;
d_mem[182] <= 13747;
d_mem[183] <= 246;
d_mem[184] <= 22461;
d_mem[185] <= 26175;
d_mem[186] <= 24195;
d_mem[187] <= 11882;
d_mem[188] <= 24021;
d_mem[189] <= 10080;
d_mem[190] <= 19856;
d_mem[191] <= 20618;
d_mem[192] <= 13930;
d_mem[193] <= 21122;
d_mem[194] <= 4097;
d_mem[195] <= 8352;
d_mem[196] <= 6986;
d_mem[197] <= 20948;
d_mem[198] <= 17277;
d_mem[199] <= 15391;
d_mem[200] <= 15049;
d_mem[201] <= 14472;
d_mem[202] <= 2631;
d_mem[203] <= 10038;
d_mem[204] <= 304;
d_mem[205] <= 5268;
d_mem[206] <= 15764;
d_mem[207] <= 13248;
d_mem[208] <= 14062;
d_mem[209] <= 26012;
d_mem[210] <= 15753;
d_mem[211] <= 9513;
d_mem[212] <= 8998;
d_mem[213] <= 23102;
d_mem[214] <= 16357;
d_mem[215] <= 4459;
d_mem[216] <= 21931;
d_mem[217] <= 992;
d_mem[218] <= 10133;
d_mem[219] <= 16993;
d_mem[220] <= 24552;
d_mem[221] <= 10716;
d_mem[222] <= 18989;
d_mem[223] <= 14251;
d_mem[224] <= 7574;
d_mem[225] <= 10984;
d_mem[226] <= 15291;
d_mem[227] <= 5347;
d_mem[228] <= 8289;
d_mem[229] <= 21285;
d_mem[230] <= 12428;
d_mem[231] <= 7685;
d_mem[232] <= 21841;
d_mem[233] <= 6240;
d_mem[234] <= 22656;
d_mem[235] <= 20171;
d_mem[236] <= 13789;
d_mem[237] <= 8641;
d_mem[238] <= 22109;
d_mem[239] <= 20576;
d_mem[240] <= 15370;
d_mem[241] <= 4228;
d_mem[242] <= 18931;
d_mem[243] <= 1807;
d_mem[244] <= 14482;
d_mem[245] <= 5946;
d_mem[246] <= 8520;
d_mem[247] <= 8452;
d_mem[248] <= 14498;
d_mem[249] <= 10773;
d_mem[250] <= 12607;
d_mem[251] <= 8331;
d_mem[252] <= 14193;
d_mem[253] <= 5027;
d_mem[254] <= 2137;
d_mem[255] <= 8767;
d_mem[256] <= 14078;
d_mem[257] <= 178;
d_mem[258] <= 22650;
d_mem[259] <= 10726;
d_mem[260] <= 5016;
d_mem[261] <= 11567;
d_mem[262] <= 4050;
d_mem[263] <= 12255;
d_mem[264] <= 15827;
d_mem[265] <= 22477;
d_mem[266] <= 20029;
d_mem[267] <= 21474;
d_mem[268] <= 4092;
d_mem[269] <= 11546;
d_mem[270] <= 9134;
d_mem[271] <= 7800;
d_mem[272] <= 1691;
d_mem[273] <= 16935;
d_mem[274] <= 17581;
d_mem[275] <= 23270;
d_mem[276] <= 10910;
d_mem[277] <= 5226;
d_mem[278] <= 5069;
d_mem[279] <= 22482;
d_mem[280] <= 9618;
d_mem[281] <= 23270;
d_mem[282] <= 2032;
d_mem[283] <= 24358;
d_mem[284] <= 8326;
d_mem[285] <= 25077;
d_mem[286] <= 3850;
d_mem[287] <= 5006;
d_mem[288] <= 1250;
d_mem[289] <= 17618;
d_mem[290] <= 8735;
d_mem[291] <= 3530;
d_mem[292] <= 9770;
d_mem[293] <= 5909;
d_mem[294] <= 25167;
d_mem[295] <= 22766;
d_mem[296] <= 914;
d_mem[297] <= 21332;
d_mem[298] <= 136;
d_mem[299] <= 14577;
d_mem[300] <= 24079;
d_mem[301] <= 15212;
d_mem[302] <= 10579;
d_mem[303] <= 18952;
d_mem[304] <= 24179;
d_mem[305] <= 162;
d_mem[306] <= 13053;
d_mem[307] <= 5027;
d_mem[308] <= 5935;
d_mem[309] <= 2589;
d_mem[310] <= 16431;
d_mem[311] <= 2967;
d_mem[312] <= 2836;
d_mem[313] <= 18916;
d_mem[314] <= 4212;
d_mem[315] <= 4423;
d_mem[316] <= 3966;
d_mem[317] <= 6056;
d_mem[318] <= 19073;
d_mem[319] <= 2510;
d_mem[320] <= 21952;
d_mem[321] <= 8709;
d_mem[322] <= 19945;
d_mem[323] <= 3923;
d_mem[324] <= 5079;
d_mem[325] <= 14908;
d_mem[326] <= 2153;
d_mem[327] <= 19840;
d_mem[328] <= 2274;
d_mem[329] <= 26128;
d_mem[330] <= 12008;
d_mem[331] <= 3262;
d_mem[332] <= 378;
d_mem[333] <= 17313;
d_mem[334] <= 17786;
d_mem[335] <= 6256;
d_mem[336] <= 12181;
d_mem[337] <= 4843;
d_mem[338] <= 9544;
d_mem[339] <= 3766;
d_mem[340] <= 21201;
d_mem[341] <= 23029;
d_mem[342] <= 13437;
d_mem[343] <= 18989;
d_mem[344] <= 2048;
d_mem[345] <= 14214;
d_mem[346] <= 9823;
d_mem[347] <= 2201;
d_mem[348] <= 6025;
d_mem[349] <= 2526;
d_mem[350] <= 9282;
d_mem[351] <= 20140;
d_mem[352] <= 18994;
d_mem[353] <= 13127;
d_mem[354] <= 21106;
d_mem[355] <= 8961;
d_mem[356] <= 16525;
d_mem[357] <= 25450;
d_mem[358] <= 26;
d_mem[359] <= 15154;
d_mem[360] <= 25072;
d_mem[361] <= 23118;
d_mem[362] <= 14219;
d_mem[363] <= 17912;
d_mem[364] <= 1654;
d_mem[365] <= 3577;
d_mem[366] <= 20507;
d_mem[367] <= 5520;
d_mem[368] <= 15291;
d_mem[369] <= 15769;
d_mem[370] <= 16935;
d_mem[371] <= 21174;
d_mem[372] <= 7454;
d_mem[373] <= 15317;
d_mem[374] <= 499;
d_mem[375] <= 13111;
d_mem[376] <= 1255;
d_mem[377] <= 12066;
d_mem[378] <= 3482;
d_mem[379] <= 24788;
d_mem[380] <= 12785;
d_mem[381] <= 12964;
d_mem[382] <= 1413;
d_mem[383] <= 20118;
d_mem[384] <= 2883;
d_mem[385] <= 1575;
d_mem[386] <= 23512;
d_mem[387] <= 4323;
d_mem[388] <= 1628;
d_mem[389] <= 18075;
d_mem[390] <= 17938;
d_mem[391] <= 7375;
d_mem[392] <= 5226;
d_mem[393] <= 20124;
d_mem[394] <= 11813;
d_mem[395] <= 1549;
d_mem[396] <= 20050;
d_mem[397] <= 20423;
d_mem[398] <= 15795;
d_mem[399] <= 22157;
d_mem[400] <= 19472;
d_mem[401] <= 18653;
d_mem[402] <= 7144;
d_mem[403] <= 12360;
d_mem[404] <= 4948;
d_mem[405] <= 15223;
d_mem[406] <= 9518;
d_mem[407] <= 8189;
d_mem[408] <= 12423;
d_mem[409] <= 25209;
d_mem[410] <= 5016;
d_mem[411] <= 15370;
d_mem[412] <= 1344;
d_mem[413] <= 23885;
d_mem[414] <= 9071;
d_mem[415] <= 13085;
d_mem[416] <= 11020;
d_mem[417] <= 9949;
d_mem[418] <= 15070;
d_mem[419] <= 16814;
d_mem[420] <= 25230;
d_mem[421] <= 2158;
d_mem[422] <= 24373;
d_mem[423] <= 23391;
d_mem[424] <= 22330;
d_mem[425] <= 25881;
d_mem[426] <= 9870;
d_mem[427] <= 14298;
d_mem[428] <= 20428;
d_mem[429] <= 11808;
d_mem[430] <= 1927;
d_mem[431] <= 4948;
d_mem[432] <= 23044;
d_mem[433] <= 9035;
d_mem[434] <= 10311;
d_mem[435] <= 26117;
d_mem[436] <= 3692;
d_mem[437] <= 11351;
d_mem[438] <= 903;
d_mem[439] <= 17334;
d_mem[440] <= 4543;
d_mem[441] <= 17587;
d_mem[442] <= 7585;
d_mem[443] <= 10800;
d_mem[444] <= 12045;
d_mem[445] <= 6539;
d_mem[446] <= 9576;
d_mem[447] <= 5547;
d_mem[448] <= 14366;
d_mem[449] <= 7989;
d_mem[450] <= 12796;
d_mem[451] <= 9329;
d_mem[452] <= 17024;
d_mem[453] <= 24342;
d_mem[454] <= 24205;
d_mem[455] <= 1092;
d_mem[456] <= 16373;
d_mem[457] <= 18164;
d_mem[458] <= 19147;
d_mem[459] <= 2668;
d_mem[460] <= 10737;
d_mem[461] <= 8651;
d_mem[462] <= 22488;
d_mem[463] <= 6413;
d_mem[464] <= 10416;
d_mem[465] <= 18564;
d_mem[466] <= 4081;
d_mem[467] <= 3703;
d_mem[468] <= 4391;
d_mem[469] <= 23969;
d_mem[470] <= 23990;
d_mem[471] <= 26086;
d_mem[472] <= 14298;
d_mem[473] <= 961;
d_mem[474] <= 1560;
d_mem[475] <= 22004;
d_mem[476] <= 8698;
d_mem[477] <= 22456;
d_mem[478] <= 25072;
d_mem[479] <= 26159;
d_mem[480] <= 13594;
d_mem[481] <= 1533;
d_mem[482] <= 24846;
d_mem[483] <= 12165;
d_mem[484] <= 7942;
d_mem[485] <= 11425;
d_mem[486] <= 8993;
d_mem[487] <= 26207;
d_mem[488] <= 3955;
d_mem[489] <= 16468;
d_mem[490] <= 15270;
d_mem[491] <= 6839;
d_mem[492] <= 6818;
d_mem[493] <= 6455;
d_mem[494] <= 17208;
d_mem[495] <= 16814;
d_mem[496] <= 7427;
d_mem[497] <= 3824;
d_mem[498] <= 840;
d_mem[499] <= 199;
d_mem[500] <= 10033;
d_mem[501] <= 23349;
d_mem[502] <= 21458;
d_mem[503] <= 15879;
d_mem[504] <= 11945;
d_mem[505] <= 11472;
d_mem[506] <= 23801;
d_mem[507] <= 25072;
d_mem[508] <= 18380;
d_mem[509] <= 12838;
d_mem[510] <= 15123;
d_mem[511] <= 3325;
d_mem[512] <= 7186;
d_mem[513] <= 23612;
d_mem[514] <= 12512;
d_mem[515] <= 6245;
d_mem[516] <= 7727;
d_mem[517] <= 6272;
d_mem[518] <= 15585;
d_mem[519] <= 11031;
d_mem[520] <= 14030;
d_mem[521] <= 23864;
d_mem[522] <= 2994;
d_mem[523] <= 14781;
d_mem[524] <= 17875;
d_mem[525] <= 17833;
d_mem[526] <= 210;
d_mem[527] <= 13368;
d_mem[528] <= 26018;
d_mem[529] <= 21763;
d_mem[530] <= 1313;
d_mem[531] <= 1160;
d_mem[532] <= 10863;
d_mem[533] <= 25976;
d_mem[534] <= 10374;
d_mem[535] <= 25456;
d_mem[536] <= 9161;
d_mem[537] <= 7401;
d_mem[538] <= 20675;
d_mem[539] <= 22692;
d_mem[540] <= 20696;
d_mem[541] <= 14797;
d_mem[542] <= 7601;
d_mem[543] <= 24531;
d_mem[544] <= 20528;
d_mem[545] <= 309;
d_mem[546] <= 15927;
d_mem[547] <= 13631;
d_mem[548] <= 16678;
d_mem[549] <= 13500;
d_mem[550] <= 14992;
d_mem[551] <= 21332;
d_mem[552] <= 14739;
d_mem[553] <= 18080;
d_mem[554] <= 16179;
d_mem[555] <= 5914;
d_mem[556] <= 20208;
d_mem[557] <= 11057;
d_mem[558] <= 19194;
d_mem[559] <= 16079;
d_mem[560] <= 14498;
d_mem[561] <= 22367;
d_mem[562] <= 20796;
d_mem[563] <= 9812;
d_mem[564] <= 11136;
d_mem[565] <= 3987;
d_mem[566] <= 6198;
d_mem[567] <= 13463;
d_mem[568] <= 18254;
d_mem[569] <= 9366;
d_mem[570] <= 8504;
d_mem[571] <= 6167;
d_mem[572] <= 3172;
d_mem[573] <= 15470;
d_mem[574] <= 23134;
d_mem[575] <= 24473;
d_mem[576] <= 840;
d_mem[577] <= 13405;
d_mem[578] <= 2101;
d_mem[579] <= 18732;
d_mem[580] <= 7816;
d_mem[581] <= 7937;
d_mem[582] <= 2878;
d_mem[583] <= 25424;
d_mem[584] <= 7222;
d_mem[585] <= 1213;
d_mem[586] <= 1050;
d_mem[587] <= 12507;
d_mem[588] <= 12549;
d_mem[589] <= 24027;
d_mem[590] <= 6282;
d_mem[591] <= 20197;
d_mem[592] <= 24053;
d_mem[593] <= 23627;
d_mem[594] <= 4270;
d_mem[595] <= 20828;
d_mem[596] <= 25802;
d_mem[597] <= 10878;
d_mem[598] <= 8262;
d_mem[599] <= 13232;
d_mem[600] <= 23092;
d_mem[601] <= 950;
d_mem[602] <= 9250;
d_mem[603] <= 25293;
d_mem[604] <= 25482;
d_mem[605] <= 10196;
d_mem[606] <= 16510;
d_mem[607] <= 24247;
d_mem[608] <= 15569;
d_mem[609] <= 11456;
d_mem[610] <= 7979;
d_mem[611] <= 9108;
d_mem[612] <= 23501;
d_mem[613] <= 4969;
d_mem[614] <= 8494;
d_mem[615] <= 13768;
d_mem[616] <= 13416;
d_mem[617] <= 23186;
d_mem[618] <= 26259;
d_mem[619] <= 14634;
d_mem[620] <= 24993;
d_mem[621] <= 6697;
d_mem[622] <= 17718;
d_mem[623] <= 11225;
d_mem[624] <= 15979;
d_mem[625] <= 12559;
d_mem[626] <= 1838;
d_mem[627] <= 11845;
d_mem[628] <= 22383;
d_mem[629] <= 12186;
d_mem[630] <= 11477;
d_mem[631] <= 24878;
d_mem[632] <= 10984;
d_mem[633] <= 25261;
d_mem[634] <= 21495;
d_mem[635] <= 7795;
d_mem[636] <= 9329;
d_mem[637] <= 11414;
d_mem[638] <= 5163;
d_mem[639] <= 5657;
d_mem[640] <= 24914;
d_mem[641] <= 11026;
d_mem[642] <= 6282;
d_mem[643] <= 10653;
d_mem[644] <= 23470;
d_mem[645] <= 13631;
d_mem[646] <= 18684;
d_mem[647] <= 25235;
d_mem[648] <= 23990;
d_mem[649] <= 6350;
d_mem[650] <= 5752;
d_mem[651] <= 12896;
d_mem[652] <= 16736;
d_mem[653] <= 22267;
d_mem[654] <= 3057;
d_mem[655] <= 25892;
d_mem[656] <= 4727;
d_mem[657] <= 3361;
d_mem[658] <= 16730;
d_mem[659] <= 7280;
d_mem[660] <= 2563;
d_mem[661] <= 7911;
d_mem[662] <= 11976;
d_mem[663] <= 6424;
d_mem[664] <= 19577;
d_mem[665] <= 21279;
d_mem[666] <= 17581;
d_mem[667] <= 6949;
d_mem[668] <= 3934;
d_mem[669] <= 25214;
d_mem[670] <= 16662;
d_mem[671] <= 19551;
d_mem[672] <= 4260;
d_mem[673] <= 9418;
d_mem[674] <= 16216;
d_mem[675] <= 2679;
d_mem[676] <= 25088;
d_mem[677] <= 10343;
d_mem[678] <= 21521;
d_mem[679] <= 1250;
d_mem[680] <= 6792;
d_mem[681] <= 14188;
d_mem[682] <= 16720;
d_mem[683] <= 5394;
d_mem[684] <= 4585;
d_mem[685] <= 16909;
d_mem[686] <= 803;
d_mem[687] <= 3472;
d_mem[688] <= 19935;
d_mem[689] <= 8347;
d_mem[690] <= 14240;
d_mem[691] <= 5620;
d_mem[692] <= 2174;
d_mem[693] <= 3435;
d_mem[694] <= 24930;
d_mem[695] <= 16830;
d_mem[696] <= 22913;
d_mem[697] <= 7711;
d_mem[698] <= 19152;
d_mem[699] <= 21038;
d_mem[700] <= 22777;
d_mem[701] <= 10537;
d_mem[702] <= 21631;
d_mem[703] <= 10416;
d_mem[704] <= 20118;
d_mem[705] <= 4874;
d_mem[706] <= 19042;
d_mem[707] <= 2847;
d_mem[708] <= 1071;
d_mem[709] <= 14902;
d_mem[710] <= 24100;
d_mem[711] <= 10427;
d_mem[712] <= 6293;
d_mem[713] <= 3262;
d_mem[714] <= 19625;
d_mem[715] <= 5116;
d_mem[716] <= 13253;
d_mem[717] <= 330;
d_mem[718] <= 9859;
d_mem[719] <= 10448;
d_mem[720] <= 7422;
d_mem[721] <= 11682;
d_mem[722] <= 3314;
d_mem[723] <= 20229;
d_mem[724] <= 21358;
d_mem[725] <= 6702;
d_mem[726] <= 11388;
d_mem[727] <= 3067;
d_mem[728] <= 7364;
d_mem[729] <= 13090;
d_mem[730] <= 7091;
d_mem[731] <= 1780;
d_mem[732] <= 11272;
d_mem[733] <= 19420;
d_mem[734] <= 829;
d_mem[735] <= 9140;
d_mem[736] <= 22866;
d_mem[737] <= 11094;
d_mem[738] <= 13410;
d_mem[739] <= 8499;
d_mem[740] <= 10847;
d_mem[741] <= 26217;
d_mem[742] <= 20203;
d_mem[743] <= 15034;
d_mem[744] <= 6135;
d_mem[745] <= 7007;
d_mem[746] <= 18579;
d_mem[747] <= 4748;
d_mem[748] <= 11089;
d_mem[749] <= 8247;
d_mem[750] <= 21910;
d_mem[751] <= 4123;
d_mem[752] <= 24347;
d_mem[753] <= 10159;
d_mem[754] <= 13116;
d_mem[755] <= 551;
d_mem[756] <= 18417;
d_mem[757] <= 7580;
d_mem[758] <= 9586;
d_mem[759] <= 1307;
d_mem[760] <= 15296;
d_mem[761] <= 11525;
d_mem[762] <= 20476;
d_mem[763] <= 18002;
d_mem[764] <= 22162;
d_mem[765] <= 24368;
d_mem[766] <= 15018;
d_mem[767] <= 1686;
d_mem[768] <= 1491;
d_mem[769] <= 19709;
d_mem[770] <= 12559;
d_mem[771] <= 26243;
d_mem[772] <= 25587;
d_mem[773] <= 22298;
d_mem[774] <= 25466;
d_mem[775] <= 5578;
d_mem[776] <= 11241;
d_mem[777] <= 21826;
d_mem[778] <= 8835;
d_mem[779] <= 9040;
d_mem[780] <= 24074;
d_mem[781] <= 20318;
d_mem[782] <= 761;
d_mem[783] <= 13663;
d_mem[784] <= 20612;
d_mem[785] <= 13248;
d_mem[786] <= 20323;
d_mem[787] <= 15969;
d_mem[788] <= 9287;
d_mem[789] <= 24773;
d_mem[790] <= 824;
d_mem[791] <= 5636;
d_mem[792] <= 5274;
d_mem[793] <= 16047;
d_mem[794] <= 25266;
d_mem[795] <= 24914;
d_mem[796] <= 13841;
d_mem[797] <= 9371;
d_mem[798] <= 12680;
d_mem[799] <= 13521;
d_mem[800] <= 24405;
d_mem[801] <= 2652;
d_mem[802] <= 11955;
d_mem[803] <= 4381;
d_mem[804] <= 12638;
d_mem[805] <= 1103;
d_mem[806] <= 13116;
d_mem[807] <= 330;
d_mem[808] <= 3708;
d_mem[809] <= 24846;
d_mem[810] <= 225;
d_mem[811] <= 25892;
d_mem[812] <= 4459;
d_mem[813] <= 18774;
d_mem[814] <= 1980;
d_mem[815] <= 26128;
d_mem[816] <= 11020;
d_mem[817] <= 25687;
d_mem[818] <= 19015;
d_mem[819] <= 22230;
d_mem[820] <= 3246;
d_mem[821] <= 6377;
d_mem[822] <= 17340;
d_mem[823] <= 367;
d_mem[824] <= 20917;
d_mem[825] <= 26065;
d_mem[826] <= 25461;
d_mem[827] <= 16042;
d_mem[828] <= 2316;
d_mem[829] <= 7422;
d_mem[830] <= 19483;
d_mem[831] <= 19562;
d_mem[832] <= 3073;
d_mem[833] <= 17660;
d_mem[834] <= 18821;
d_mem[835] <= 22892;
d_mem[836] <= 14314;
d_mem[837] <= 15653;
d_mem[838] <= 7317;
d_mem[839] <= 22372;
d_mem[840] <= 18789;
d_mem[841] <= 23218;
d_mem[842] <= 11078;
d_mem[843] <= 25555;
d_mem[844] <= 20287;
d_mem[845] <= 5757;
d_mem[846] <= 9639;
d_mem[847] <= 12722;
d_mem[848] <= 13799;
d_mem[849] <= 3435;
d_mem[850] <= 20660;
d_mem[851] <= 13410;
d_mem[852] <= 5762;
d_mem[853] <= 8121;
d_mem[854] <= 19877;
d_mem[855] <= 9339;
d_mem[856] <= 10322;
d_mem[857] <= 12838;
d_mem[858] <= 7270;
d_mem[859] <= 5415;
d_mem[860] <= 26049;
d_mem[861] <= 4354;
d_mem[862] <= 6986;
d_mem[863] <= 7947;
d_mem[864] <= 7159;
d_mem[865] <= 18338;
d_mem[866] <= 8068;
d_mem[867] <= 4491;
d_mem[868] <= 22677;
d_mem[869] <= 7585;
d_mem[870] <= 1560;
d_mem[871] <= 14671;
d_mem[872] <= 25314;
d_mem[873] <= 19373;
d_mem[874] <= 18947;
d_mem[875] <= 4869;
d_mem[876] <= 13353;
d_mem[877] <= 15049;
d_mem[878] <= 6203;
d_mem[879] <= 1985;
d_mem[880] <= 18742;
d_mem[881] <= 2810;
d_mem[882] <= 1602;
d_mem[883] <= 13001;
d_mem[884] <= 12838;
d_mem[885] <= 3398;
d_mem[886] <= 11209;
d_mem[887] <= 23176;
d_mem[888] <= 15564;
d_mem[889] <= 24521;
d_mem[890] <= 9481;
d_mem[891] <= 1786;
d_mem[892] <= 23507;
d_mem[893] <= 14839;
d_mem[894] <= 6582;
d_mem[895] <= 709;
d_mem[896] <= 13642;
d_mem[897] <= 20665;
d_mem[898] <= 10001;
d_mem[899] <= 9182;
d_mem[900] <= 25960;
d_mem[901] <= 17235;
d_mem[902] <= 2269;
d_mem[903] <= 18322;
d_mem[904] <= 18984;
d_mem[905] <= 2132;
d_mem[906] <= 21610;
d_mem[907] <= 19183;
d_mem[908] <= 9329;
d_mem[909] <= 18753;
d_mem[910] <= 10553;
d_mem[911] <= 6613;
d_mem[912] <= 4543;
d_mem[913] <= 2253;
d_mem[914] <= 19824;
d_mem[915] <= 21384;
d_mem[916] <= 4943;
d_mem[917] <= 17891;
d_mem[918] <= 24878;
d_mem[919] <= 4937;
d_mem[920] <= 535;
d_mem[921] <= 16867;
d_mem[922] <= 577;
d_mem[923] <= 10947;
d_mem[924] <= 17051;
d_mem[925] <= 20933;
d_mem[926] <= 24605;
d_mem[927] <= 12922;
d_mem[928] <= 120;
d_mem[929] <= 15259;
d_mem[930] <= 5242;
d_mem[931] <= 1171;
d_mem[932] <= 20297;
d_mem[933] <= 23260;
d_mem[934] <= 11462;
d_mem[935] <= 17786;
d_mem[936] <= 10689;
d_mem[937] <= 25508;
d_mem[938] <= 5147;
d_mem[939] <= 4580;
d_mem[940] <= 18348;
d_mem[941] <= 8882;
d_mem[942] <= 25419;
d_mem[943] <= 23444;
d_mem[944] <= 241;
d_mem[945] <= 1759;
d_mem[946] <= 4869;
d_mem[947] <= 1276;
d_mem[948] <= 17324;
d_mem[949] <= 9492;
d_mem[950] <= 2290;
d_mem[951] <= 12990;
d_mem[952] <= 5752;
d_mem[953] <= 10805;
d_mem[954] <= 13342;
d_mem[955] <= 7138;
d_mem[956] <= 1765;
d_mem[957] <= 24605;
d_mem[958] <= 7653;
d_mem[959] <= 20392;
d_mem[960] <= 173;
d_mem[961] <= 17124;
d_mem[962] <= 6356;
d_mem[963] <= 5962;
d_mem[964] <= 6907;
d_mem[965] <= 6870;
d_mem[966] <= 12207;
d_mem[967] <= 19656;
d_mem[968] <= 20854;
d_mem[969] <= 10269;
d_mem[970] <= 25587;
d_mem[971] <= 19898;
d_mem[972] <= 3099;
d_mem[973] <= 6277;
d_mem[974] <= 22845;
d_mem[975] <= 1596;
d_mem[976] <= 330;
d_mem[977] <= 5074;
d_mem[978] <= 23244;
d_mem[979] <= 20807;
d_mem[980] <= 5442;
d_mem[981] <= 89;
d_mem[982] <= 14608;
d_mem[983] <= 2169;
d_mem[984] <= 10915;
d_mem[985] <= 25366;
d_mem[986] <= 7427;
d_mem[987] <= 23097;
d_mem[988] <= 12985;
d_mem[989] <= 18674;
d_mem[990] <= 8593;
d_mem[991] <= 3692;
d_mem[992] <= 4381;
d_mem[993] <= 1386;
d_mem[994] <= 25949;
d_mem[995] <= 8593;
d_mem[996] <= 21174;
d_mem[997] <= 12827;
d_mem[998] <= 15044;
d_mem[999] <= 147;
d_mem[1000] <= 9092;
d_mem[1001] <= 21190;
d_mem[1002] <= 13295;
d_mem[1003] <= 16420;
d_mem[1004] <= 10133;
d_mem[1005] <= 16525;
d_mem[1006] <= 2379;
d_mem[1007] <= 8473;
d_mem[1008] <= 8840;
d_mem[1009] <= 11225;
d_mem[1010] <= 24741;
d_mem[1011] <= 19914;
d_mem[1012] <= 20355;
d_mem[1013] <= 25403;
d_mem[1014] <= 23491;
d_mem[1015] <= 8063;
d_mem[1016] <= 5263;
d_mem[1017] <= 10632;
d_mem[1018] <= 698;
d_mem[1019] <= 15916;
d_mem[1020] <= 20801;
d_mem[1021] <= 13053;
d_mem[1022] <= 23339;
d_mem[1023] <= 18096;
d_mem[1024] <= 18506;//*/
  
  /*/64badde
  d_mem[0] <= 16'hfffe;
  d_mem[1] <= 16'hfffe;
  d_mem[2] <= 16'hfffe;
  d_mem[3] <= 16'h0000;
  d_mem[4] <= 16'hffff;
  d_mem[5] <= 16'hffff;
  d_mem[6] <= 16'hffff;
  d_mem[7] <= 16'h0000;//*/
  //*/init_test
  /*d_mem[0] <= 16'hfffd;
  d_mem[1] <= 16'h0004;
  d_mem[2] <= 16'h0005;
  d_mem[3] <= 16'hc369;
  d_mem[4] <= 16'h69c3;
  d_mem[5] <= 16'h0041;
  d_mem[6] <= 16'hffff;
  d_mem[7] <= 16'h0001;//*/
  end
  else
  begin
    if(dwe) d_mem[addr] <= wdata;
	 else 
		 begin 
		 rdata <= d_mem[addr]; 
		 tocache <= {d_mem[{addr[15:2],2'b00}],d_mem[{addr[15:2],2'b01}],d_mem[{addr[15:2],2'b10}],d_mem[{addr[15:2],2'b11}]};
		 end
  end
end

endmodule
